module INV_VERILOG(PSW0, LED0);
    input  PSW0;
    output LED0;

    assign LED0 = ~PSW0;

endmodule
